// ----  Probes  ----
`define PROBE_ADDR      pd1.addr
`define PROBE_DATA_IN   pd1.data_in
`define PROBE_DATA_OUT  pd1.data_out
`define PROBE_READ_EN   pd1.read_en
`define PROBE_WRITE_EN  pd1.write_en

`define PROBE_F_PC      pd1.fetch_pc
`define PROBE_F_INSN    pd1.fetch_insn
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd1
// ----  Top module  ----
